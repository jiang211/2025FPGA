module fft_top #(
    parameter integer DATAIN_WIDTH    = 16   ,                           
    parameter integer DATAOUT_WIDTH   = 32   ,                           
    parameter integer USER_WIDTH      = 16                           
)
(
    input                      clk                            ,
    input                      rst_n                          ,
 
    // �ⲿ���ݽӿ�      
    input                      data_input_start_flag          ,   //fft_modulus_fifo�洢���������־
    input                      wd_en                          ,   //fft ipдʹ��
    input  [DATAIN_WIDTH-1:0]  wd_data                        ,   //д�ź�����
    output                     rd_en                          ,   //��ʹ��
    output [DATAOUT_WIDTH-1:0] fft_amplitude_frequency_data       //�����Ƶ����

   );

wire                          xn_axi4s_data_tvalid         ;
wire   [DATAIN_WIDTH*2-1:0]   xn_axi4s_data_tdata          ;
wire                          xn_axi4s_data_tlast          ;
wire                          xn_axi4s_data_tready         ;
wire                          xn_axi4s_cfg_tvalid          ;
wire                          xn_axi4s_cfg_tdata           ;
wire                          xk_axi4s_data_tvalid         ;
wire   [DATAOUT_WIDTH*2-1:0]  xk_axi4s_data_tdata          ;
wire                          xk_axi4s_data_tlast          ;
wire   [USER_WIDTH-1:0]       xk_axi4s_data_tuser          ;
wire   [2:0]                  alm                          ;
wire                          stat                         ;
                                                           
wire  [DATAOUT_WIDTH-1:0]     out_fft_data_re              ;
wire  [DATAOUT_WIDTH-1:0]     out_fft_data_im              ;
wire                          source_valid                 ;

wire                          source_sop                   ;
wire                          source_eop                   ;


fft_axi_master #(
    .DATAIN_WIDTH        (DATAIN_WIDTH        ),                           
    .DATAOUT_WIDTH       (DATAOUT_WIDTH       ),                           
    .USER_WIDTH          (USER_WIDTH          )                        
)
u_fft_axi_master
(
    .clk                 (clk                 ),
    .rst_n               (rst_n               ),                      
    .wd_en               (wd_en               ),   //дʹ��
    .rd_en               (source_valid        ),   //��ʹ��
    .wd_data             (wd_data             ),   //д�ź�����   
    .out_fft_data_re     (out_fft_data_re     ),   //���fft���ݣ�ʵ����
    .out_fft_data_im     (out_fft_data_im     ),   //���fft���ݣ��鲿��
    .fft_sop             (source_sop          ),
    .fft_eop             (source_eop          ),

    .i_axi4s_data_tvalid (xn_axi4s_data_tvalid),
    .i_axi4s_data_tdata  (xn_axi4s_data_tdata ),
    .i_axi4s_data_tlast  (xn_axi4s_data_tlast ),
    .o_axi4s_data_tready (xn_axi4s_data_tready),
    .i_axi4s_cfg_tvalid  (xn_axi4s_cfg_tvalid ),
    .i_axi4s_cfg_tdata   (xn_axi4s_cfg_tdata  ),
                        
    .o_axi4s_data_tvalid (xk_axi4s_data_tvalid),
    .o_axi4s_data_tdata  (xk_axi4s_data_tdata ),
    .o_axi4s_data_tlast  (xk_axi4s_data_tlast ),
    .o_axi4s_data_tuser  (xk_axi4s_data_tuser ),
    .o_alm               (alm                 ),
    .o_stat              (stat                )

   );


fft_data_modulus u_fft_data_modulus(
    .clk                    (clk                          ),
    .rst_n                  (rst_n                        ),
    //FFT ST�ӿ�          
    .source_real            (out_fft_data_re              ),
    .source_imag            (out_fft_data_im              ),
    .source_sop             (source_sop                   ),
    .source_eop             (source_eop                   ),
    .source_valid           (source_valid                 ),
    //ȡģ���������ݽӿ�        
    .data_modulus           (fft_amplitude_frequency_data ),  
    .data_modulus_valid     (rd_en                        ),
    //�û��ӿ�
    .data_input_start_flag  (data_input_start_flag        )
   );


fft_demo_00  u_fft_wrapper ( 
    .i_aclk                 (clk                 ),

    .i_axi4s_data_tvalid    (xn_axi4s_data_tvalid),
    .i_axi4s_data_tdata     (xn_axi4s_data_tdata ),
    .i_axi4s_data_tlast     (xn_axi4s_data_tlast ),
    .o_axi4s_data_tready    (xn_axi4s_data_tready),
    .i_axi4s_cfg_tvalid     (xn_axi4s_cfg_tvalid ),
    .i_axi4s_cfg_tdata      (xn_axi4s_cfg_tdata  ),
    .o_axi4s_data_tvalid    (xk_axi4s_data_tvalid),
    .o_axi4s_data_tdata     (xk_axi4s_data_tdata ),
    .o_axi4s_data_tlast     (xk_axi4s_data_tlast ),
    .o_axi4s_data_tuser     (xk_axi4s_data_tuser ),
    .o_alm                  (alm                 ),
    .o_stat                 (stat                )
);



endmodule