module sin_lut #(
    parameter DATA_WIDTH = 8
) (
    input  [DATA_WIDTH:0] addr,
    output reg [DATA_WIDTH-1:0] data
);

always @(*) begin
    case (addr)
0 : data = 8'h80;
1 : data = 8'h81;
2 : data = 8'h83;
3 : data = 8'h84;
4 : data = 8'h86;
5 : data = 8'h87;
6 : data = 8'h89;
7 : data = 8'h8A;
8 : data = 8'h8C;
9 : data = 8'h8E;
10 : data = 8'h8F;
11 : data = 8'h91;
12 : data = 8'h92;
13 : data = 8'h94;
14 : data = 8'h95;
15 : data = 8'h97;
16 : data = 8'h98;
17 : data = 8'h9A;
18 : data = 8'h9C;
19 : data = 8'h9D;
20 : data = 8'h9F;
21 : data = 8'hA0;
22 : data = 8'hA2;
23 : data = 8'hA3;
24 : data = 8'hA5;
25 : data = 8'hA6;
26 : data = 8'hA8;
27 : data = 8'hA9;
28 : data = 8'hAB;
29 : data = 8'hAC;
30 : data = 8'hAE;
31 : data = 8'hAF;
32 : data = 8'hB0;
33 : data = 8'hB2;
34 : data = 8'hB3;
35 : data = 8'hB5;
36 : data = 8'hB6;
37 : data = 8'hB8;
38 : data = 8'hB9;
39 : data = 8'hBA;
40 : data = 8'hBC;
41 : data = 8'hBD;
42 : data = 8'hBF;
43 : data = 8'hC0;
44 : data = 8'hC1;
45 : data = 8'hC3;
46 : data = 8'hC4;
47 : data = 8'hC5;
48 : data = 8'hC7;
49 : data = 8'hC8;
50 : data = 8'hC9;
51 : data = 8'hCA;
52 : data = 8'hCC;
53 : data = 8'hCD;
54 : data = 8'hCE;
55 : data = 8'hCF;
56 : data = 8'hD1;
57 : data = 8'hD2;
58 : data = 8'hD3;
59 : data = 8'hD4;
60 : data = 8'hD5;
61 : data = 8'hD7;
62 : data = 8'hD8;
63 : data = 8'hD9;
64 : data = 8'hDA;
65 : data = 8'hDB;
66 : data = 8'hDC;
67 : data = 8'hDD;
68 : data = 8'hDE;
69 : data = 8'hDF;
70 : data = 8'hE0;
71 : data = 8'hE1;
72 : data = 8'hE2;
73 : data = 8'hE3;
74 : data = 8'hE4;
75 : data = 8'hE5;
76 : data = 8'hE6;
77 : data = 8'hE7;
78 : data = 8'hE8;
79 : data = 8'hE9;
80 : data = 8'hEA;
81 : data = 8'hEB;
82 : data = 8'hEC;
83 : data = 8'hEC;
84 : data = 8'hED;
85 : data = 8'hEE;
86 : data = 8'hEF;
87 : data = 8'hF0;
88 : data = 8'hF0;
89 : data = 8'hF1;
90 : data = 8'hF2;
91 : data = 8'hF3;
92 : data = 8'hF3;
93 : data = 8'hF4;
94 : data = 8'hF5;
95 : data = 8'hF5;
96 : data = 8'hF6;
97 : data = 8'hF6;
98 : data = 8'hF7;
99 : data = 8'hF7;
100 : data = 8'hF8;
101 : data = 8'hF9;
102 : data = 8'hF9;
103 : data = 8'hFA;
104 : data = 8'hFA;
105 : data = 8'hFA;
106 : data = 8'hFB;
107 : data = 8'hFB;
108 : data = 8'hFC;
109 : data = 8'hFC;
110 : data = 8'hFC;
111 : data = 8'hFD;
112 : data = 8'hFD;
113 : data = 8'hFD;
114 : data = 8'hFE;
115 : data = 8'hFE;
116 : data = 8'hFE;
117 : data = 8'hFE;
118 : data = 8'hFF;
119 : data = 8'hFF;
120 : data = 8'hFF;
121 : data = 8'hFF;
122 : data = 8'hFF;
123 : data = 8'hFF;
124 : data = 8'hFF;
125 : data = 8'hFF;
126 : data = 8'hFF;
127 : data = 8'hFF;
128 : data = 8'hFF;
129 : data = 8'hFF;
130 : data = 8'hFF;
131 : data = 8'hFF;
132 : data = 8'hFF;
133 : data = 8'hFF;
134 : data = 8'hFF;
135 : data = 8'hFF;
136 : data = 8'hFF;
137 : data = 8'hFF;
138 : data = 8'hFF;
139 : data = 8'hFE;
140 : data = 8'hFE;
141 : data = 8'hFE;
142 : data = 8'hFE;
143 : data = 8'hFD;
144 : data = 8'hFD;
145 : data = 8'hFD;
146 : data = 8'hFC;
147 : data = 8'hFC;
148 : data = 8'hFC;
149 : data = 8'hFB;
150 : data = 8'hFB;
151 : data = 8'hFA;
152 : data = 8'hFA;
153 : data = 8'hFA;
154 : data = 8'hF9;
155 : data = 8'hF9;
156 : data = 8'hF8;
157 : data = 8'hF7;
158 : data = 8'hF7;
159 : data = 8'hF6;
160 : data = 8'hF6;
161 : data = 8'hF5;
162 : data = 8'hF5;
163 : data = 8'hF4;
164 : data = 8'hF3;
165 : data = 8'hF3;
166 : data = 8'hF2;
167 : data = 8'hF1;
168 : data = 8'hF0;
169 : data = 8'hF0;
170 : data = 8'hEF;
171 : data = 8'hEE;
172 : data = 8'hED;
173 : data = 8'hEC;
174 : data = 8'hEC;
175 : data = 8'hEB;
176 : data = 8'hEA;
177 : data = 8'hE9;
178 : data = 8'hE8;
179 : data = 8'hE7;
180 : data = 8'hE6;
181 : data = 8'hE5;
182 : data = 8'hE4;
183 : data = 8'hE3;
184 : data = 8'hE2;
185 : data = 8'hE1;
186 : data = 8'hE0;
187 : data = 8'hDF;
188 : data = 8'hDE;
189 : data = 8'hDD;
190 : data = 8'hDC;
191 : data = 8'hDB;
192 : data = 8'hDA;
193 : data = 8'hD9;
194 : data = 8'hD8;
195 : data = 8'hD7;
196 : data = 8'hD5;
197 : data = 8'hD4;
198 : data = 8'hD3;
199 : data = 8'hD2;
200 : data = 8'hD1;
201 : data = 8'hCF;
202 : data = 8'hCE;
203 : data = 8'hCD;
204 : data = 8'hCC;
205 : data = 8'hCA;
206 : data = 8'hC9;
207 : data = 8'hC8;
208 : data = 8'hC7;
209 : data = 8'hC5;
210 : data = 8'hC4;
211 : data = 8'hC3;
212 : data = 8'hC1;
213 : data = 8'hC0;
214 : data = 8'hBF;
215 : data = 8'hBD;
216 : data = 8'hBC;
217 : data = 8'hBA;
218 : data = 8'hB9;
219 : data = 8'hB8;
220 : data = 8'hB6;
221 : data = 8'hB5;
222 : data = 8'hB3;
223 : data = 8'hB2;
224 : data = 8'hB0;
225 : data = 8'hAF;
226 : data = 8'hAE;
227 : data = 8'hAC;
228 : data = 8'hAB;
229 : data = 8'hA9;
230 : data = 8'hA8;
231 : data = 8'hA6;
232 : data = 8'hA5;
233 : data = 8'hA3;
234 : data = 8'hA2;
235 : data = 8'hA0;
236 : data = 8'h9F;
237 : data = 8'h9D;
238 : data = 8'h9C;
239 : data = 8'h9A;
240 : data = 8'h98;
241 : data = 8'h97;
242 : data = 8'h95;
243 : data = 8'h94;
244 : data = 8'h92;
245 : data = 8'h91;
246 : data = 8'h8F;
247 : data = 8'h8E;
248 : data = 8'h8C;
249 : data = 8'h8A;
250 : data = 8'h89;
251 : data = 8'h87;
252 : data = 8'h86;
253 : data = 8'h84;
254 : data = 8'h83;
255 : data = 8'h81;
256 : data = 8'h80;
257 : data = 8'h7E;
258 : data = 8'h7C;
259 : data = 8'h7B;
260 : data = 8'h79;
261 : data = 8'h78;
262 : data = 8'h76;
263 : data = 8'h75;
264 : data = 8'h73;
265 : data = 8'h71;
266 : data = 8'h70;
267 : data = 8'h6E;
268 : data = 8'h6D;
269 : data = 8'h6B;
270 : data = 8'h6A;
271 : data = 8'h68;
272 : data = 8'h67;
273 : data = 8'h65;
274 : data = 8'h63;
275 : data = 8'h62;
276 : data = 8'h60;
277 : data = 8'h5F;
278 : data = 8'h5D;
279 : data = 8'h5C;
280 : data = 8'h5A;
281 : data = 8'h59;
282 : data = 8'h57;
283 : data = 8'h56;
284 : data = 8'h54;
285 : data = 8'h53;
286 : data = 8'h51;
287 : data = 8'h50;
288 : data = 8'h4F;
289 : data = 8'h4D;
290 : data = 8'h4C;
291 : data = 8'h4A;
292 : data = 8'h49;
293 : data = 8'h47;
294 : data = 8'h46;
295 : data = 8'h45;
296 : data = 8'h43;
297 : data = 8'h42;
298 : data = 8'h40;
299 : data = 8'h3F;
300 : data = 8'h3E;
301 : data = 8'h3C;
302 : data = 8'h3B;
303 : data = 8'h3A;
304 : data = 8'h38;
305 : data = 8'h37;
306 : data = 8'h36;
307 : data = 8'h35;
308 : data = 8'h33;
309 : data = 8'h32;
310 : data = 8'h31;
311 : data = 8'h30;
312 : data = 8'h2E;
313 : data = 8'h2D;
314 : data = 8'h2C;
315 : data = 8'h2B;
316 : data = 8'h2A;
317 : data = 8'h28;
318 : data = 8'h27;
319 : data = 8'h26;
320 : data = 8'h25;
321 : data = 8'h24;
322 : data = 8'h23;
323 : data = 8'h22;
324 : data = 8'h21;
325 : data = 8'h20;
326 : data = 8'h1F;
327 : data = 8'h1E;
328 : data = 8'h1D;
329 : data = 8'h1C;
330 : data = 8'h1B;
331 : data = 8'h1A;
332 : data = 8'h19;
333 : data = 8'h18;
334 : data = 8'h17;
335 : data = 8'h16;
336 : data = 8'h15;
337 : data = 8'h14;
338 : data = 8'h13;
339 : data = 8'h13;
340 : data = 8'h12;
341 : data = 8'h11;
342 : data = 8'h10;
343 : data = 8'h0F;
344 : data = 8'h0F;
345 : data = 8'h0E;
346 : data = 8'h0D;
347 : data = 8'h0C;
348 : data = 8'h0C;
349 : data = 8'h0B;
350 : data = 8'h0A;
351 : data = 8'h0A;
352 : data = 8'h09;
353 : data = 8'h09;
354 : data = 8'h08;
355 : data = 8'h08;
356 : data = 8'h07;
357 : data = 8'h06;
358 : data = 8'h06;
359 : data = 8'h05;
360 : data = 8'h05;
361 : data = 8'h05;
362 : data = 8'h04;
363 : data = 8'h04;
364 : data = 8'h03;
365 : data = 8'h03;
366 : data = 8'h03;
367 : data = 8'h02;
368 : data = 8'h02;
369 : data = 8'h02;
370 : data = 8'h01;
371 : data = 8'h01;
372 : data = 8'h01;
373 : data = 8'h01;
374 : data = 8'h00;
375 : data = 8'h00;
376 : data = 8'h00;
377 : data = 8'h00;
378 : data = 8'h00;
379 : data = 8'h00;
380 : data = 8'h00;
381 : data = 8'h00;
382 : data = 8'h00;
383 : data = 8'h00;
384 : data = 8'h00;
385 : data = 8'h00;
386 : data = 8'h00;
387 : data = 8'h00;
388 : data = 8'h00;
389 : data = 8'h00;
390 : data = 8'h00;
391 : data = 8'h00;
392 : data = 8'h00;
393 : data = 8'h00;
394 : data = 8'h00;
395 : data = 8'h01;
396 : data = 8'h01;
397 : data = 8'h01;
398 : data = 8'h01;
399 : data = 8'h02;
400 : data = 8'h02;
401 : data = 8'h02;
402 : data = 8'h03;
403 : data = 8'h03;
404 : data = 8'h03;
405 : data = 8'h04;
406 : data = 8'h04;
407 : data = 8'h05;
408 : data = 8'h05;
409 : data = 8'h05;
410 : data = 8'h06;
411 : data = 8'h06;
412 : data = 8'h07;
413 : data = 8'h08;
414 : data = 8'h08;
415 : data = 8'h09;
416 : data = 8'h09;
417 : data = 8'h0A;
418 : data = 8'h0A;
419 : data = 8'h0B;
420 : data = 8'h0C;
421 : data = 8'h0C;
422 : data = 8'h0D;
423 : data = 8'h0E;
424 : data = 8'h0F;
425 : data = 8'h0F;
426 : data = 8'h10;
427 : data = 8'h11;
428 : data = 8'h12;
429 : data = 8'h13;
430 : data = 8'h13;
431 : data = 8'h14;
432 : data = 8'h15;
433 : data = 8'h16;
434 : data = 8'h17;
435 : data = 8'h18;
436 : data = 8'h19;
437 : data = 8'h1A;
438 : data = 8'h1B;
439 : data = 8'h1C;
440 : data = 8'h1D;
441 : data = 8'h1E;
442 : data = 8'h1F;
443 : data = 8'h20;
444 : data = 8'h21;
445 : data = 8'h22;
446 : data = 8'h23;
447 : data = 8'h24;
448 : data = 8'h25;
449 : data = 8'h26;
450 : data = 8'h27;
451 : data = 8'h28;
452 : data = 8'h2A;
453 : data = 8'h2B;
454 : data = 8'h2C;
455 : data = 8'h2D;
456 : data = 8'h2E;
457 : data = 8'h30;
458 : data = 8'h31;
459 : data = 8'h32;
460 : data = 8'h33;
461 : data = 8'h35;
462 : data = 8'h36;
463 : data = 8'h37;
464 : data = 8'h38;
465 : data = 8'h3A;
466 : data = 8'h3B;
467 : data = 8'h3C;
468 : data = 8'h3E;
469 : data = 8'h3F;
470 : data = 8'h40;
471 : data = 8'h42;
472 : data = 8'h43;
473 : data = 8'h45;
474 : data = 8'h46;
475 : data = 8'h47;
476 : data = 8'h49;
477 : data = 8'h4A;
478 : data = 8'h4C;
479 : data = 8'h4D;
480 : data = 8'h4F;
481 : data = 8'h50;
482 : data = 8'h51;
483 : data = 8'h53;
484 : data = 8'h54;
485 : data = 8'h56;
486 : data = 8'h57;
487 : data = 8'h59;
488 : data = 8'h5A;
489 : data = 8'h5C;
490 : data = 8'h5D;
491 : data = 8'h5F;
492 : data = 8'h60;
493 : data = 8'h62;
494 : data = 8'h63;
495 : data = 8'h65;
496 : data = 8'h67;
497 : data = 8'h68;
498 : data = 8'h6A;
499 : data = 8'h6B;
500 : data = 8'h6D;
501 : data = 8'h6E;
502 : data = 8'h70;
503 : data = 8'h71;
504 : data = 8'h73;
505 : data = 8'h75;
506 : data = 8'h76;
507 : data = 8'h78;
508 : data = 8'h79;
509 : data = 8'h7B;
510 : data = 8'h7C;
511 : data = 8'h7E;
        default: data = 8'h00;
    endcase
end

endmodule
