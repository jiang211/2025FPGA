module top #(
    parameter PH_W = 32,
    parameter DT_W = 8
) (
    input  wire                clk,
    input  wire                rst_n,
    
    input  wire [PH_W-1:0]     freq_word,
    input  wire [DT_W-1:0]     amplitude,  // 峰值（正数）
    input gate,

    input [DT_W -1 : 0] wave_in,
    output [1:0] wave_type
);
localparam SAD_FREQ = 97656; 

localparam THRESHOLD = 10;

localparam IDLE = 0;
localparam START_MATCHING = 1;
localparam FINISH_MATCHING = 2;

//gate 开启之后开始寻找峰值
reg [1:0] matching_gate;
reg [7:0] cycle_cnt;
always @(posedge clk) begin
    if(!gate)begin
        matching_gate <= IDLE;
        cycle_cnt <= 0;
    end else begin
        case (matching_gate)
            IDLE :begin
             if(wave_in - amplitude <= THRESHOLD || amplitude - wave_in <= THRESHOLD) matching_gate <= START_MATCHING;
            end 
            START_MATCHING : begin

             cycle_cnt <= cycle_cnt + 1;
             if(cycle_cnt == 255) matching_gate <= FINISH_MATCHING;   

            end
            FINISH_MATCHING : begin

            end
            default: matching_gate <= IDLE;
        endcase
    end
end

//从输入波形的峰值开始进行模板匹配
reg [7:0] wave_reg0;
reg [7:0] wave_reg1;
reg [7:0] wave_reg2;
always @(posedge clk) begin
    wave_reg0 <= wave_in;
    wave_reg1 <= wave_reg0;
    wave_reg2 <= wave_reg1;
end


//对输入波形进行求导
wire [7:0] dwave;
divirative u_dut (
    .clk_50M        (clk),
    .rst_n      (matching_gate),

    .valid      (matching_gate),
    .wave_data  (wave_in),
    .fifo_dout  (dwave),

    .circle_cnt (circle_cnt),
    .output_valid(output_valid)
);

//产生一个三角波模板
wire [7:0] tri_wave;
wire [7:0] tri_wave_270;
wire [7:0] sqr_wave;
wire [7:0] dsqr_wave;

triangle_dds dut0 (
    .clk(clk),
    .rst_n(matching_gate),

    .freq_word(freq_word),
    .amplitude(amplitude),
    .wave_out(tri_wave),
    .wave_out_270(tri_wave_270)

);

//产生方波模板
sqr_wave_gen dut1 (
    .clk(clk),
    .rst_n(matching_gate),
    
    .freq_word(freq_word),
    .amplitude(amplitude),
    .sel_phase(0),
    .wave_out(sqr_wave)
);

//产生三角波的求导波


sqr_wave_gen dut2 (
    .clk(clk),
    .rst_n(matching_gate),
    
    .freq_word(freq_word),
    .amplitude(freq_word/SAD_FREQ +128),
    .sel_phase(0),
    .wave_out(dsqr_wave)
);
//模板匹配
template_match u_template_match (
    .clk        (clk),
    .rst_n      (rst_n),

    .wave_valid (matching_gate),
    .type_valid (type_valid),

    .tri_template (tri_wave),
    .sqr_template (sqr_wave),
    .sin_template (tri_wave),
    .dtri_template (dsqr_wave),
    .dsin_template (tri_wave_270),

    .wave_in    (wave_reg2),
    .dwave_in   (dwave),
    .wave_type  (wave_type)
);


endmodule