module tri_lut #(
    parameter DATA_WIDTH = 8
) (
    input  [DATA_WIDTH-1:0] addr,
    output [DATA_WIDTH-1:0] data
);

always @(*) begin
    case (addr)
0 : data = 0
1 : data = 1
2 : data = 2
3 : data = 3
4 : data = 4
5 : data = 5
6 : data = 6
7 : data = 7
8 : data = 8
9 : data = 9
10 : data = 10
11 : data = 11
12 : data = 12
13 : data = 13
14 : data = 14
15 : data = 15
16 : data = 16
17 : data = 17
18 : data = 18
19 : data = 19
20 : data = 20
21 : data = 21
22 : data = 22
23 : data = 23
24 : data = 24
25 : data = 25
26 : data = 26
27 : data = 27
28 : data = 28
29 : data = 29
30 : data = 30
31 : data = 31
32 : data = 32
33 : data = 33
34 : data = 34
35 : data = 35
36 : data = 36
37 : data = 37
38 : data = 38
39 : data = 39
40 : data = 40
41 : data = 41
42 : data = 42
43 : data = 43
44 : data = 44
45 : data = 45
46 : data = 46
47 : data = 47
48 : data = 48
49 : data = 49
50 : data = 50
51 : data = 51
52 : data = 52
53 : data = 53
54 : data = 54
55 : data = 55
56 : data = 56
57 : data = 57
58 : data = 58
59 : data = 59
60 : data = 60
61 : data = 61
62 : data = 62
63 : data = 63
64 : data = 64
65 : data = 65
66 : data = 66
67 : data = 67
68 : data = 68
69 : data = 69
70 : data = 70
71 : data = 71
72 : data = 72
73 : data = 73
74 : data = 74
75 : data = 75
76 : data = 76
77 : data = 77
78 : data = 78
79 : data = 79
80 : data = 80
81 : data = 81
82 : data = 82
83 : data = 83
84 : data = 84
85 : data = 85
86 : data = 86
87 : data = 87
88 : data = 88
89 : data = 89
90 : data = 90
91 : data = 91
92 : data = 92
93 : data = 93
94 : data = 94
95 : data = 95
96 : data = 96
97 : data = 97
98 : data = 98
99 : data = 99
100 : data = 100
101 : data = 101
102 : data = 102
103 : data = 103
104 : data = 104
105 : data = 105
106 : data = 106
107 : data = 107
108 : data = 108
109 : data = 109
110 : data = 110
111 : data = 111
112 : data = 112
113 : data = 113
114 : data = 114
115 : data = 115
116 : data = 116
117 : data = 117
118 : data = 118
119 : data = 119
120 : data = 120
121 : data = 121
122 : data = 122
123 : data = 123
124 : data = 124
125 : data = 125
126 : data = 126
127 : data = 127
128 : data = 128
129 : data = 129
130 : data = 130
131 : data = 131
132 : data = 132
133 : data = 133
134 : data = 134
135 : data = 135
136 : data = 136
137 : data = 137
138 : data = 138
139 : data = 139
140 : data = 140
141 : data = 141
142 : data = 142
143 : data = 143
144 : data = 144
145 : data = 145
146 : data = 146
147 : data = 147
148 : data = 148
149 : data = 149
150 : data = 150
151 : data = 151
152 : data = 152
153 : data = 153
154 : data = 154
155 : data = 155
156 : data = 156
157 : data = 157
158 : data = 158
159 : data = 159
160 : data = 160
161 : data = 161
162 : data = 162
163 : data = 163
164 : data = 164
165 : data = 165
166 : data = 166
167 : data = 167
168 : data = 168
169 : data = 169
170 : data = 170
171 : data = 171
172 : data = 172
173 : data = 173
174 : data = 174
175 : data = 175
176 : data = 176
177 : data = 177
178 : data = 178
179 : data = 179
180 : data = 180
181 : data = 181
182 : data = 182
183 : data = 183
184 : data = 184
185 : data = 185
186 : data = 186
187 : data = 187
188 : data = 188
189 : data = 189
190 : data = 190
191 : data = 191
192 : data = 192
193 : data = 193
194 : data = 194
195 : data = 195
196 : data = 196
197 : data = 197
198 : data = 198
199 : data = 199
200 : data = 200
201 : data = 201
202 : data = 202
203 : data = 203
204 : data = 204
205 : data = 205
206 : data = 206
207 : data = 207
208 : data = 208
209 : data = 209
210 : data = 210
211 : data = 211
212 : data = 212
213 : data = 213
214 : data = 214
215 : data = 215
216 : data = 216
217 : data = 217
218 : data = 218
219 : data = 219
220 : data = 220
221 : data = 221
222 : data = 222
223 : data = 223
224 : data = 224
225 : data = 225
226 : data = 226
227 : data = 227
228 : data = 228
229 : data = 229
230 : data = 230
231 : data = 231
232 : data = 232
233 : data = 233
234 : data = 234
235 : data = 235
236 : data = 236
237 : data = 237
238 : data = 238
239 : data = 239
240 : data = 240
241 : data = 241
242 : data = 242
243 : data = 243
244 : data = 244
245 : data = 245
246 : data = 246
247 : data = 247
248 : data = 248
249 : data = 249
250 : data = 250
251 : data = 251
252 : data = 252
253 : data = 253
254 : data = 254
257 : data = 255
258 : data = 254
259 : data = 253
260 : data = 252
261 : data = 251
262 : data = 250
263 : data = 249
264 : data = 248
265 : data = 247
266 : data = 246
267 : data = 245
268 : data = 244
269 : data = 243
270 : data = 242
271 : data = 241
272 : data = 240
273 : data = 239
274 : data = 238
275 : data = 237
276 : data = 236
277 : data = 235
278 : data = 234
279 : data = 233
280 : data = 232
281 : data = 231
282 : data = 230
283 : data = 229
284 : data = 228
285 : data = 227
286 : data = 226
287 : data = 225
288 : data = 224
289 : data = 223
290 : data = 222
291 : data = 221
292 : data = 220
293 : data = 219
294 : data = 218
295 : data = 217
296 : data = 216
297 : data = 215
298 : data = 214
299 : data = 213
300 : data = 212
301 : data = 211
302 : data = 210
303 : data = 209
304 : data = 208
305 : data = 207
306 : data = 206
307 : data = 205
308 : data = 204
309 : data = 203
310 : data = 202
311 : data = 201
312 : data = 200
313 : data = 199
314 : data = 198
315 : data = 197
316 : data = 196
317 : data = 195
318 : data = 194
319 : data = 193
320 : data = 192
321 : data = 191
322 : data = 190
323 : data = 189
324 : data = 188
325 : data = 187
326 : data = 186
327 : data = 185
328 : data = 184
329 : data = 183
330 : data = 182
331 : data = 181
332 : data = 180
333 : data = 179
334 : data = 178
335 : data = 177
336 : data = 176
337 : data = 175
338 : data = 174
339 : data = 173
340 : data = 172
341 : data = 171
342 : data = 170
343 : data = 169
344 : data = 168
345 : data = 167
346 : data = 166
347 : data = 165
348 : data = 164
349 : data = 163
350 : data = 162
351 : data = 161
352 : data = 160
353 : data = 159
354 : data = 158
355 : data = 157
356 : data = 156
357 : data = 155
358 : data = 154
359 : data = 153
360 : data = 152
361 : data = 151
362 : data = 150
363 : data = 149
364 : data = 148
365 : data = 147
366 : data = 146
367 : data = 145
368 : data = 144
369 : data = 143
370 : data = 142
371 : data = 141
372 : data = 140
373 : data = 139
374 : data = 138
375 : data = 137
376 : data = 136
377 : data = 135
378 : data = 134
379 : data = 133
380 : data = 132
381 : data = 131
382 : data = 130
383 : data = 129
384 : data = 128
385 : data = 127
386 : data = 126
387 : data = 125
388 : data = 124
389 : data = 123
390 : data = 122
391 : data = 121
392 : data = 120
393 : data = 119
394 : data = 118
395 : data = 117
396 : data = 116
397 : data = 115
398 : data = 114
399 : data = 113
400 : data = 112
401 : data = 111
402 : data = 110
403 : data = 109
404 : data = 108
405 : data = 107
406 : data = 106
407 : data = 105
408 : data = 104
409 : data = 103
410 : data = 102
411 : data = 101
412 : data = 100
413 : data = 99
414 : data = 98
415 : data = 97
416 : data = 96
417 : data = 95
418 : data = 94
419 : data = 93
420 : data = 92
421 : data = 91
422 : data = 90
423 : data = 89
424 : data = 88
425 : data = 87
426 : data = 86
427 : data = 85
428 : data = 84
429 : data = 83
430 : data = 82
431 : data = 81
432 : data = 80
433 : data = 79
434 : data = 78
435 : data = 77
436 : data = 76
437 : data = 75
438 : data = 74
439 : data = 73
440 : data = 72
441 : data = 71
442 : data = 70
443 : data = 69
444 : data = 68
445 : data = 67
446 : data = 66
447 : data = 65
448 : data = 64
449 : data = 63
450 : data = 62
451 : data = 61
452 : data = 60
453 : data = 59
454 : data = 58
455 : data = 57
456 : data = 56
457 : data = 55
458 : data = 54
459 : data = 53
460 : data = 52
461 : data = 51
462 : data = 50
463 : data = 49
464 : data = 48
465 : data = 47
466 : data = 46
467 : data = 45
468 : data = 44
469 : data = 43
470 : data = 42
471 : data = 41
472 : data = 40
473 : data = 39
474 : data = 38
475 : data = 37
476 : data = 36
477 : data = 35
478 : data = 34
479 : data = 33
480 : data = 32
481 : data = 31
482 : data = 30
483 : data = 29
484 : data = 28
485 : data = 27
486 : data = 26
487 : data = 25
488 : data = 24
489 : data = 23
490 : data = 22
491 : data = 21
492 : data = 20
493 : data = 19
494 : data = 18
495 : data = 17
496 : data = 16
497 : data = 15
498 : data = 14
499 : data = 13
500 : data = 12
501 : data = 11
502 : data = 10
503 : data = 9
504 : data = 8
505 : data = 7
506 : data = 6
507 : data = 5
508 : data = 4
509 : data = 3
510 : data = 2
511 : data = 1
512 : data = 0
        default: data = 8'h00;
    endcase
end

endmodule
